// save_settings.v

module hamnn
