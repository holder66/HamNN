// multiple_test.v
module hamnn

// test_multiple_classifiers 
fn test_multiple_classifiers() {
	
}