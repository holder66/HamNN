// load_file_test.v
module hamnn

// test_load_instances_file 
fn test_load_instances_file() ? {
	
}