// oxplot.v

module hamnn

