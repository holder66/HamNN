// oxplot.v

module hamnn