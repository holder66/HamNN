// multiple.v

module hamnn