// save.v
module tools

// import os
