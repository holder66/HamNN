// display_test.v
module display
