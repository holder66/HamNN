// multiple.v

module hamnn

// multiple_classifier_classify
fn multiple_classifier_classify(classifiers []Classifier, instances [][]u8, opts Options) ClassifyResult {
	mut mcr := ClassifyResult{}
	return mcr
}
