// display_test.v
module display

// test_display 
fn test_display() {
	
}