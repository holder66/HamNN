// append_test.v
module append
