// display.v
module display

import tools
// import os

// display
pub fn display(opts tools.Options) {
}
