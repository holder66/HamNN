// plot_test.v
module tools

// test_two_array_sort
fn test_two_array_sort() {
	two_array_sort([1., 2, 3], [4., 5, 6])
}