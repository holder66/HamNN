// append.v
module append

import tools

// append 
pub fn append(cl tools.Classifier, opts tools.Options) ?tools.Classifier {
	return cl
}